//拿AI写了一个imem用于测试功能
module imem (
    input  logic [31:0] addr,
    output logic [31:0] instr
);

    logic [31:0] mem [0:255];

    initial begin
        integer i;
        for (i = 0; i < 256; i = i + 1)
            mem[i] = 32'b0;

        // =========================
        // 初始化数据区（dmem[0] = 5）
        // =========================
        // lw  $t0, 0($zero)
        mem[0] = 32'b100011_00000_01000_0000000000000000;

        // =========================
        // load-use hazard（必须 stall）
        // =========================
        // add $t1, $t0, $t0   -> 10
        mem[1] = 32'b000000_01000_01000_01001_00000_100000;

        // =========================
        // forwarding（不用 stall）
        // =========================
        // add $t2, $t0, $t0   -> 10
        mem[2] = 32'b000000_01000_01000_01010_00000_100000;

        // =========================
        // addi
        // =========================
        // addi $t3, $zero, 3
        mem[3] = 32'b001000_00000_01011_0000000000000011;

        // =========================
        // andi / ori / xor
        // =========================
        // andi $t4, $t3, 1   -> 1
        mem[4] = 32'b001100_01011_01100_0000000000000001;

        // ori  $t5, $t3, 2   -> 3
        mem[5] = 32'b001101_01011_01101_0000000000000010;

        // xor  $t6, $t4, $t5 -> 1 ^ 3 = 2
        mem[6] = 32'b000000_01100_01101_01110_00000_100110;

        // =========================
        // lui
        // =========================
        // lui $t7, 0x1234 -> 0x12340000
        mem[7] = 32'b001111_00000_01111_0001001000110100;

        // =========================
        // slt
        // =========================
        // slt $s0, $t4, $t5  (1 < 3) -> 1
        mem[8] = 32'b000000_01100_01101_10000_00000_101010;

        // =========================
        // beq taken（触发 flush）
        // =========================
        // beq $s0, $t4, +1   (1 == 1) -> taken
        mem[9]  = 32'b000100_10000_01100_0000000000000001;

        // ❌ 这条应被 flush
        // addi $s1, $zero, 99
        mem[10] = 32'b001000_00000_10001_0000000001100011;

        // =========================
        // 正常继续
        // =========================
        // addi $s1, $zero, 7
        mem[11] = 32'b001000_00000_10001_0000000000000111;

        // =========================
        // sw / lw
        // =========================
        // sw $s1, 4($zero)
        mem[12] = 32'b101011_00000_10001_0000000000000100;

        // lw $s2, 4($zero)
        mem[13] = 32'b100011_00000_10010_0000000000000100;
    end

    assign instr = mem[addr[9:2]];

endmodule
